module programCounterAdder(
    input [3:0] I,
    output [3:0] O
);
    assign O = I + 1;
endmodule